
// 4 OP | 12 Immediate

localparam OP_NOP   = 0;
localparam OP_CLEAR = 1;

localparam OP_POS   = 12;
localparam OP_SIZE  = 4;
